// Code your design here
`include "mc_top.v"